library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_arith.all;

entity if_id_reg is port
(
	CLK		: in std_logic;
   PC_if		: in std_logic_vector(31 downto 0);
	INST_if	: in std_logic_vector(31 downto 0);
   PC_id		: out std_logic_vector(31 downto 0);
	INST_id	: out std_logic_vector(31 downto 0)
);
end if_id_reg;

architecture behavior of if_id_reg is
begin
	process(CLK)
	begin
		if CLK'event and CLK = '1' then
			PC_id <= PC_if;
			INST_id <= INST_if;
		end if;
	end process;
end behavior;
